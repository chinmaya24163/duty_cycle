\TLV_version 1d: tl-x.org
\SV
/* verilator lint_off UNUSED*/  /* verilator lint_off DECLFILENAME*/  /* verilator lint_off BLKSEQ*/  /* verilator lint_off WIDTH*/  /* verilator lint_off SELRANGE*/  /* verilator lint_off PINCONNECTEMPTY*/  /* verilator lint_off DEFPARAM*/  /* verilator lint_off IMPLICIT*/  /* verilator lint_off COMBDLY*/  /* verilator lint_off SYNCASYNCNET*/  /* verilator lint_off UNOPTFLAT */  /* verilator lint_off UNSIGNED*/  /* verilator lint_off CASEINCOMPLETE*/  /* verilator lint_off UNDRIVEN*/  /* verilator lint_off VARHIDDEN*/  /* verilator lint_off CASEX*/  /* verilator lint_off CASEOVERLAP*/  /* verilator lint_off PINMISSING*/  /* verilator lint_off LATCH*/  /* verilator lint_off BLKANDNBLK*/  /* verilator lint_off MULTIDRIVEN*/  /* verilator lint_off NULLPORT*/  /* verilator lint_off EOFNEWLINE*/  /* verilator lint_off WIDTHCONCAT*/  /* verilator lint_off ASSIGNDLY*/  /* verilator lint_off MODDUP*/  /* verilator lint_off STMTDLY*/  /* verilator lint_off LITENDIAN*/  /* verilator lint_off INITIALDLY*/  

//Your Verilog/System Verilog Code Starts Here:
`timescale 1ns / 1ps

module duty_cycle(input clk, output reg out);
    reg [1:0] curr_state = 0; 
    reg [1:0] next_state;

    always @(posedge clk) begin
        curr_state <= next_state;
    end

    always @(*) begin
        case(curr_state)
            2'b00: out = 1;
            2'b01: out = 0;
            2'b10: out = 0;
            2'b11: out = 0;
            default: out = 0;
        endcase
    end

    always @(*) begin
        next_state = curr_state + 1;
    end    
endmodule

//Top Module Code Starts here:
	module top(input logic clk, input logic reset, input logic [31:0] cyc_cnt, output logic passed, output logic failed);
//The $random() can be replaced if user wants to assign values
		logic out_sig;

		duty_cycle duty_cycle_inst(
			.clk(clk),
			.out(out_sig)
		);

		always_ff @(posedge clk) begin
			if (reset) begin
				passed <= 0;
				failed <= 0;
			end else begin
				if (cyc_cnt > 20) begin
					passed <= 1;
					failed <= 0;
				end
			end
		end
	endmodule